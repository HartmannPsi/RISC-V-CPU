`inlcude "../macros.v"

module ReservationStation();
endmodule